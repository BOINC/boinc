#Swedish language.ini file

#pay attention to the NOTE in the [MENU- ] section

#PROJECT_ID
[HEADER-Projects]
Title=Projekt
Project=Projekt
Account=Konto
Total Credit=Total Arbete
Avg. Credit=Genomsnittligt Arbete
Resource Share=Resurs

#RESULT_ID
[HEADER-Work]
Title=Arbete
Project=Projekt
Application=Program
Name=Namn
CPU time=CPU Tid
Progress=Utf�rt
To Completion=Till Klar
Status=Status

#XFER_ID
[HEADER-Transfers]
Title=�verf�ringar
Project=Projekt
File=Fil
Progress=Utf�rt
Size=Storlek
Time=Tid
Speed=Hastighet
Status=Status

#MESSAGE_ID
[HEADER-Messages]
Title=Meddelanden
Project=Projekt
Time=Tid
Message=Besked

#USAGE_ID
[HEADER-Disk]
Title=Disk
Free space: not available for use=Ledig Storlek: Kan Ej Anv�ndas
Free space: available for use=Ledig Storlek: Kan Anv�ndas
Used space: other than BOINC=Anv�nd Storlek: Ut�ver BOINC
Used space: BOINC=Anv�nd Storlek: BOINC
Used space:=Anv�nd Storlek

#miscellaneous text
[HEADER-MISC]
New=Ny
Running=K�r
Ready to run=Klar
Computation done=Ber�kningar Utf�rt
Results uploaded=Resultat Skickat
Acknowledged=Bekr�ftat
Error: invalid state=Fel: Ogiltigt Tillst�nd
Completed=Utf�rt
Uploading=Laddar Upp
Downloading=Laddar Ner
Retry in=F�rs�k Igen Om
Upload failed=Uppladdning Misslyckad
Download failed=Nerladdning Misslyckad

#menu items
# NOTE: add an & (ampersand) to the letter to be used as mnemonic
#       i.e. Show Graphics=Show &Graphics
#                               ^^ the "G" will trigger the menu item
#       you can compare it with a saved language.ini.XX file
[MENU-File]
Title=&Titel
Show Graphics=&Visa Grafik
Clear Messages=Radera &Meddelanden
Clear Inactive=Radera &Inaktiva
Suspend=&Paus
Resume=&Forts�tt
Exit=&Exit

[MENU-Settings]
Title=&Inst�llningar
Login to Project...=Logga &In
Quit Project...=Logga &Ut
Proxy Server...=&Proxy

[MENU-Connection]
Title=&Anslut
Connect Now=&Anslut Nu
Hangup Connection if Dialed=&L�gg P� Vid Samtal
Confirm Before Connecting=&Bekr�fta F�re Anslutning

[MENU-Work]
Show Graphics=Visa &Grafik

[MENU-Help]
Title=&Hj�lp
About...=&Om...

[MENU-StatusIcon]
Suspend=&Paus
Resume=&Forts�tt
Exit=&Avsluta

[MENU-Project]
Relogin...=&Logga In Igen
Quit Project...=&Avsluta Projekt

[DIALOG-LOGIN]
Title=Logga In P� Projektet
URL:=Adress
Account Key:=Anv�ndar ID
OK=OK
Cancel=Avbryt
The URL for the website of the project.=Adressen Till Projektets Hemsida
The authorization code recieved in your confirmation email.=Din S�kerhetskod Som Du F�tt Via Epost

[DIALOG-QUIT]
Title=Avsluta Project
URL:=URL
Account Key:=Anv�ndar ID
OK=OK
Cancel=Avbryt
Select the project you wish to quit.=Markera Det Projekt Du Vill Avsluta

[DIALOG-CONNECT]
Title=Anslut Till N�tverket
BOINC needs to connect to the network.  May it do so now?=BOINC Beh�ver Ansluta Sig Till N�tverket.  �r Det OK Att G�ra Det ?
Don't ask this again (connect automatically)=Fr�ga Inte Fler G�nger (Anslut Automatiskt)
OK=OK
Cancel=Avbryt

[DIALOG-ABOUT]
Title=Boinc Beta Version
Berkeley Open Infrastructure for Network Computing=Berkeley Open Infrastructure for Network Computing
Open Beta=�ppen Beta-Version
OK=OK

[DIALOG-PROXY]
Title=Proxy Server Inst�llningar
Some organizations use an "HTTP proxy" or a "SOCKS proxy" (or both) for increased security.  If you need to use a proxy, fill in the information below.  If you need help, ask your System Administrator or Internet Service Provider.=Vissa Organisationer Anv�nder "HTTP Proxy" Eller "SOCKS Proxy" (Eller B�gge) F�r �kad S�kerhet. Om Du Beh�ver Anv�nda En Proxy, Fyll I Uppgifterna Nedan.  Om Du Beh�ver Hj�lp, Fr�ga Din System-Administrat�r Eller Din Internet leverant�r
HTTP Proxy=HTTP Proxy
Connect via HTTP Proxy Server=Anslut Via HTTP Proxy Server
http://=http://
Port Number:=Portnummer
SOCKS Proxy=SOCKS Proxy
Connect via SOCKS Proxy Server=Anslut Via SOCKS Proxy Server
SOCKS Host:=SOCKS V�rd
Port Number:=Portnummner
Leave these blank if not needed=L�mna Blank Om Det Inte Beh�vs
SOCKS User Name:=SOCKS Anv�ndarnamn
SOCKS Password:=SOCKS L�senord
OK=OK
Cancel=Avbryt

